//akgjagjag
