//akgjagjag
//fasgag
